`timescale 1ns/1ps

module Flush(
    input branch,
    output reg flush
);
    initial
    begin 
        flush = 1'b0;
    end
    always @(*)
    begin
      if (branch == 1'b1)
        flush = 1'b1;
      else
        flush = 1'b0;
    end

endmodule
